package enum_pkg;
  typedef enum logic [3:0] {
    Add,
    Sub,
    Leftshift,
    RightshiftArith,
    RightshiftLogic,
    And,
    Or,
    Xor,
    Equal
  } Opcode;
endpackage
