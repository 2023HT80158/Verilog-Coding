//two input AND gate

module and2 (
  	input wire A, 
  	input wire B,
  	output wire Y
);
  
	assign Y = A & B;
    
endmodule