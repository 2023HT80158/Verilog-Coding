module SRAM_tb();
  reg clk;
  reg [7:0] data_in;
  reg wr;
  reg rd;
  reg [2:0] addr;
  wire [7:0] data_out;
  
  SRAM1 dut( .clk(clk), .data_in(data_in), .wr(wr), .rd(rd), .addr(addr), .data_out(data_out));
  
  initial begin
    
   clk = 0;
  end
  always #5 clk = ~clk;
  
  initial begin
    wr = 1;
    rd = 0;
    addr = 3'b001;
    data_in = 8'b00;
    #5
    wr = 1;
    rd = 0;
    addr = 3'b001;
    data_in = 8'b00111110;
    #5
     wr = 0;
    rd = 1;
    addr = 3'b001;
    data_in = 8'b00;
   	#100  $finish ;
    
  end
  
  initial begin 
    $monitor("time = %t, wr = %d, rd = %d, data_out = %b", $time, wr, rd, data_out);
  end
endmodule
